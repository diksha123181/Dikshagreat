<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-28.4,-85.2,104.95,-153.15</PageViewport>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>38.5,-18.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>25.5,-16.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>25.5,-21.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>48.5,-18.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>22,-15.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>21.5,-20.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>55,-18</position>
<gparam>LABEL_TEXT Y=A.B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>34.5,-11.5</position>
<gparam>LABEL_TEXT AND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AE_OR2</type>
<position>39,-36.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>27,-34.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>27,-38.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>47,-36.5</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>31.5,-30.5</position>
<gparam>LABEL_TEXT OR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>22.5,-34</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>23,-38</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>55,-36</position>
<gparam>LABEL_TEXT Y= A+B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_INVERTER</type>
<position>32,-51.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>25,-51.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>40,-51.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>20.5,-51.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>44,-51</position>
<gparam>LABEL_TEXT A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>31.5,-46.5</position>
<gparam>LABEL_TEXT NOT GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>BA_NAND2</type>
<position>32,-68</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>20.5,-66.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>20.5,-69.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>41,-68</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>32,-62.5</position>
<gparam>LABEL_TEXT NAND GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>17.5,-65.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>17.5,-69.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>49,-67.5</position>
<gparam>LABEL_TEXT Y=(A.B)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>BE_NOR2</type>
<position>32,-84</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>20,-81.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>20,-86.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>41.5,-84</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>31,-78</position>
<gparam>LABEL_TEXT NOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>17,-81</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>17,-85.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>50,-83.5</position>
<gparam>LABEL_TEXT Y=(A+B)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AI_XOR2</type>
<position>31.5,-100</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>20,-97</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>20,-103</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>40.5,-100</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>31,-94</position>
<gparam>LABEL_TEXT EX-OR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>17.5,-96.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>17,-102.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>49,-99.5</position>
<gparam>LABEL_TEXT Y=A(+)B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AO_XNOR2</type>
<position>31.5,-115.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>20.5,-113</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>20.5,-118</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>GA_LED</type>
<position>39,-115.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>31.5,-109.5</position>
<gparam>LABEL_TEXT EX-NOR GATE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>17,-112.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>17,-117</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>50.5,-115</position>
<gparam>LABEL_TEXT Y=(A(+)B)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-17.5,31.5,-16.5</points>
<intersection>-17.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-17.5,35.5,-17.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-16.5,31.5,-16.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-21.5,31.5,-19.5</points>
<intersection>-21.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-19.5,35.5,-19.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-21.5,31.5,-21.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-18.5,47.5,-18.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-35.5,32.5,-34.5</points>
<intersection>-35.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-35.5,36,-35.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-34.5,32.5,-34.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-38.5,32.5,-37.5</points>
<intersection>-38.5 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-37.5,36,-37.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29,-38.5,32.5,-38.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42,-36.5,46,-36.5</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<connection>
<GID>15</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-51.5,29,-51.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-51.5,39,-51.5</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-67,25.5,-66.5</points>
<intersection>-67 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-67,29,-67</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-66.5,25.5,-66.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-69.5,25.5,-69</points>
<intersection>-69.5 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-69,29,-69</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-69.5,25.5,-69.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-68,40,-68</points>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<connection>
<GID>36</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-83,25.5,-81.5</points>
<intersection>-83 1</intersection>
<intersection>-81.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-83,29,-83</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-81.5,25.5,-81.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-86.5,25.5,-85</points>
<intersection>-86.5 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-85,29,-85</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-86.5,25.5,-86.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-84,40.5,-84</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>48</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-99,25,-97</points>
<intersection>-99 1</intersection>
<intersection>-97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-99,28.5,-99</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-97,25,-97</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-103,25,-101</points>
<intersection>-103 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-101,28.5,-101</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-103,25,-103</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-100,39.5,-100</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-114.5,25.5,-113</points>
<intersection>-114.5 1</intersection>
<intersection>-113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-114.5,28.5,-114.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-113,25.5,-113</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-118,25.5,-116.5</points>
<intersection>-118 2</intersection>
<intersection>-116.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-116.5,28.5,-116.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-118,25.5,-118</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-115.5,38,-115.5</points>
<connection>
<GID>78</GID>
<name>N_in0</name></connection>
<connection>
<GID>72</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 1>
<page 2>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 2>
<page 3>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 3>
<page 4>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 4>
<page 5>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 5>
<page 6>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 6>
<page 7>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 7>
<page 8>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 8>
<page 9>
<PageViewport>0,0,177.8,-90.6</PageViewport></page 9></circuit>